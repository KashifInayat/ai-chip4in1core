// SPDX-FileCopyrightText: 2020 Efabless Corporation
//
// Licensed under the Apache License, Version 2.0 (the "License");
// you may not use this file except in compliance with the License.
// You may obtain a copy of the License at
//
//      http://www.apache.org/licenses/LICENSE-2.0
//
// Unless required by applicable law or agreed to in writing, software
// distributed under the License is distributed on an "AS IS" BASIS,
// WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
// See the License for the specific language governing permissions and
// limitations under the License.
// SPDX-License-Identifier: Apache-2.0

`default_nettype none
/*
 *-------------------------------------------------------------
 *
 * user_project_wrapper
 *
 * This wrapper enumerates all of the pins available to the
 * user for the user project.
 *
 * An example user project is provided in this wrapper.  The
 * example should be removed and replaced with the actual
 * user project.
 *
 *-------------------------------------------------------------
 */

module user_project_wrapper #(
    parameter BITS = 32
) (
`ifdef USE_POWER_PINS
    inout vdda1,	// User area 1 3.3V supply
    inout vdda2,	// User area 2 3.3V supply
    inout vssa1,	// User area 1 analog ground
    inout vssa2,	// User area 2 analog ground
    inout vccd1,	// User area 1 1.8V supply
    inout vccd2,	// User area 2 1.8v supply
    inout vssd1,	// User area 1 digital ground
    inout vssd2,	// User area 2 digital ground
`endif

    // Wishbone Slave ports (WB MI A)
    input wb_clk_i,
    input wb_rst_i,
    input wbs_stb_i,
    input wbs_cyc_i,
    input wbs_we_i,
    input [3:0] wbs_sel_i,
    input [31:0] wbs_dat_i,
    input [31:0] wbs_adr_i,
    output wbs_ack_o,
    output [31:0] wbs_dat_o,

    // Logic Analyzer Signals
    input  [127:0] la_data_in,
    output [127:0] la_data_out,
    input  [127:0] la_oenb,

    // IOs
    input  [`MPRJ_IO_PADS-1:0] io_in,
    output [`MPRJ_IO_PADS-1:0] io_out,
    output [`MPRJ_IO_PADS-1:0] io_oeb,

    // Analog (direct connection to GPIO pad---use with caution)
    // Note that analog I/O is not available on the 7 lowest-numbered
    // GPIO pads, and so the analog_io indexing is offset from the
    // GPIO indexing by 7 (also upper 2 GPIOs do not have analog_io).
    inout [`MPRJ_IO_PADS-10:0] analog_io,

    // Independent clock (on independent integer divider)
    input   user_clock2,

    // User maskable interrupt signals
    output [2:0] user_irq
);

/*--------------------------------------*/
/* User project is instantiated  here   */
/*--------------------------------------*/

/*--------------------------------------*/
/* User project is instantiated  here   */
/*--------------------------------------*/





    FFPMAC ffpmac_0(
	    .A(la_data_in[15:0]),
	    .B(la_data_in[31:16]), 
	    .C(la_data_in[63:32]),
	    .rnd(la_oenb[1:0]),
	    .clk(clk_50),
	    .rst(wb_rst_i),
	    .result(la_data_out[31:0]));

    CLA_16 cla16_0( 
	    .OPA(la_data_in[79:64]),
	    .OPB(la_data_in[95:80]),
	    .CIN(la_oenb[2]), .PHI(la_oenb[3]),
	    .SUM_FINAL(la_data_out[47:32]),
	    .COUT_FINAL(la_data_out[48]),
	    .CLK(wb_clk_i));

    sa_2D sa2d_0( 
	

	    .AA(la_data_in[103:96]), 
	    .BB(la_data_in[111:104]), 
	    .CLK(wb_clk_i), 
	    .SHIFTEN(la_oenb[5:4]),
	    .RST(wb_rst_i), 
	    .Y(la_data_out[80:49]));

   r8_mb8 r8_mb8_0(
   
	    .mx(la_data_in[119:112]),
	    .my(la_data_in[127:120]),
	    .CLK(wb_clk_i), 
	    .RST(wb_rst_i),
	    .product_final(la_data_out[106:81]));





endmodule	// user_project_wrapper


`default_nettype wire
